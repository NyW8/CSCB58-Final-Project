module display(mode, colour, size);
	input mode, colour, size;
endmodule