module display(mode, colour, size);

endmodule