module movement(position, overlap_colour, temp);

endmodule

