module controller ();


endmodule

module setColour();

endmodule

module setSize();

endmodule

module setMode();

endmodule