module paint(SW, KEY, LEDR, HEX0, HEX1, HEX2, HEX3);
	input [17:0] SW;
	input [4:0] KEY;
	output [17:0] LEDR;
	output [6:0] HEX0;
	output [6:0] HEX1;
	output [6:0] HEX2;
	output [6:0] HEX3;
	
	/*
	This is a top-level module, please don't add code here except for testing!
	*/
endmodule